library verilog;
use verilog.vl_types.all;
entity testbench_div_hd is
end testbench_div_hd;
